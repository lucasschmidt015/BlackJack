library ieee;
use ieee.std_logic_1164.all;

entity round is
    port(
        
        clock: in std_logic;

    );
end round;

architecture behaviour of round is
begin
    process()
    begin
        
    end process;
end behaviour;