library ieee;
use ieee.std_logic_1164.all;

entity blackJack is 
    port(
        
    );
end blackJack;

architecture behaviour of blackJack is 
begin
    process()
        

    end process;
end behaviour;